// sdram.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module sdram (
		input  wire [23:0] avalon_sdram_address,       // avalon_sdram.address
		input  wire [1:0]  avalon_sdram_byteenable_n,  //             .byteenable_n
		input  wire        avalon_sdram_chipselect,    //             .chipselect
		input  wire [15:0] avalon_sdram_writedata,     //             .writedata
		input  wire        avalon_sdram_read_n,        //             .read_n
		input  wire        avalon_sdram_write_n,       //             .write_n
		output wire [15:0] avalon_sdram_readdata,      //             .readdata
		output wire        avalon_sdram_readdatavalid, //             .readdatavalid
		output wire        avalon_sdram_waitrequest,   //             .waitrequest
		input  wire        clk_clk,                    //          clk.clk
		input  wire        reset_reset_n,              //        reset.reset_n
		output wire [12:0] sdram_addr,                 //        sdram.addr
		output wire [1:0]  sdram_ba,                   //             .ba
		output wire        sdram_cas_n,                //             .cas_n
		output wire        sdram_cke,                  //             .cke
		output wire        sdram_cs_n,                 //             .cs_n
		inout  wire [15:0] sdram_dq,                   //             .dq
		output wire [1:0]  sdram_dqm,                  //             .dqm
		output wire        sdram_ras_n,                //             .ras_n
		output wire        sdram_we_n,                 //             .we_n
		input  wire        sdram_rst_reset_n           //    sdram_rst.reset_n
	);

	sdram_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (clk_clk),                    //   clk.clk
		.reset_n        (sdram_rst_reset_n),          // reset.reset_n
		.az_addr        (avalon_sdram_address),       //    s1.address
		.az_be_n        (avalon_sdram_byteenable_n),  //      .byteenable_n
		.az_cs          (avalon_sdram_chipselect),    //      .chipselect
		.az_data        (avalon_sdram_writedata),     //      .writedata
		.az_rd_n        (avalon_sdram_read_n),        //      .read_n
		.az_wr_n        (avalon_sdram_write_n),       //      .write_n
		.za_data        (avalon_sdram_readdata),      //      .readdata
		.za_valid       (avalon_sdram_readdatavalid), //      .readdatavalid
		.za_waitrequest (avalon_sdram_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                 //  wire.export
		.zs_ba          (sdram_ba),                   //      .export
		.zs_cas_n       (sdram_cas_n),                //      .export
		.zs_cke         (sdram_cke),                  //      .export
		.zs_cs_n        (sdram_cs_n),                 //      .export
		.zs_dq          (sdram_dq),                   //      .export
		.zs_dqm         (sdram_dqm),                  //      .export
		.zs_ras_n       (sdram_ras_n),                //      .export
		.zs_we_n        (sdram_we_n)                  //      .export
	);

endmodule
